* Basic Test Circuit

V1 N001 0 AC(1 0)
V2 N002 N001 1
R1 N002 N003 1k
D1 N003 N004 D
C1 N004 0 1u
R2 N004 0 100k

.ac dec 20 10 1k
.end