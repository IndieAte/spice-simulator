* Test Circuit

V1 N001 0 10
V2 N004 2
R1 N001 N002 0 10
R2 N003 0 10
NMOS N002 N004 N003

.ac dec 5 1 20
.end