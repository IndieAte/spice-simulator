* Basic Test Circuit

I1 0 N001 0.1
R1 N001 0 100
R2 N001 N002 200
D1 N002 N003 D
R3 N003 0 50

.ac dec 20 10 1k
.end