* Basic Test Circuit

V1 N001 0 5
L1 N001 N002 1m
R1 N004 0 1k
C1 N003 N004 1u
R2 N002 N003 2k
D1 N003 N005 D
D2 0 N005 D
R3 N005 0 10k

.ac dec 20 10 1k
.end