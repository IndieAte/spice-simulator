* Basic Test Circuit

V1 N001 0 10
Q1 N002 N002 N001 PNP
Q2 N003 N002 N001 PNP
R1 N002 0 9300
Q3 N003 N004 N005 NPN
R2 N003 N004 200k
R3 N005 0 1k
C1 N004 N006 1u
V2 N006 0 AC(1 0)

.ac dec 200 10 100k
.end
