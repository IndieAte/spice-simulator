* Test Circuit

* 5V -> N014
* -5V -> N015
* -IN -> N016
* OUT -> N017

Q1 N011 N016 N006 mPNP
Q2 N008 0 N006 mPNP
V2 N014 0 5
V3 0 N015 5
Q3 N006 N004 N002 mPNP
Q4 N002 N002 N014 mPNP
Q5 N004 N002 N014 mPNP
R1 N004 N015 8.6k
Q6 N008 N011 N015 mNPN
Q7 N011 N011 N015 mNPN
Q8 N003 N003 N014 mPNP
Q9 N001 N003 N014 mPNP
R4 N003 N015 9.3k
Q10 N009 N013 N015 mNPN
Q11 N009 N008 N013 mNPN
R5 N013 N015 1.5k
Q12 N014 N001 N005 mNPN
Q13 N015 N009 N010 mPNP
Q14 N001 N001 N012 mNPN
Q15 N009 N009 N012 mPNP
Q16 N009 N010 N017 mPNP
Q17 N001 N005 N017 mNPN
R9 N005 N017 2
R10 N017 N010 2
V1 N007 0 AC(10m 0)
R2 N016 N007 10k
R3 N017 N016 100k
C1 N009 N008 470p

.model mNPN NPN(Is=0.01p Bf=200 Br=1 Vaf=120 Var=120 Cjc=8p Cje=25p Fc=0.7)
.model mPNP PNP(Is=0.01p Bf=200 Br=1 Vaf=120 Var=120 Cjc=8p Cje=30p Fc=0.7)

.ac dec 100 100 10Meg
.end