* Basic Test Circuit

I1 N001 0 AC(2 45)
D1 N001 N002 1u
Q1 N002 0 1m
R1 N002 0 1k

.ac dec 20 10 1k
.end