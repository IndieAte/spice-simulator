* Test Circuit

V1 N002 0 1
V2 N001 N002 2
R1 N003 0 1
R2 N001 N003 2

.ac dec 5 1 20
.end