* Basic Test Circuit

V1 N001 0 AC(2 90)
C1 N001 N002 1u
R1 N002 0 1k
.ac dec 10 1 100

.end