* Test Circuit

V1 N001 0 50
R1 N001 N002 10k
Q1 N002 N003 0 NPN
I1 0 N003 15u

.ac dec 5 1 20
.end