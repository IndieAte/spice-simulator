* Basic Test Circuit

V1 0 N001 5
R1 N001 N002 5k
R2 N002 N003 200k
V2 N004 0 AC(0.1 0)
C1 N004 N003 1u
Q1 N002 N003 N005 PNP
R3 N005 0 1k

.ac dec 20 10 10k
.end
