* Basic Test Circuit

v1 0 N001 AC(1 180)
R1 N001 N002 1
R2 N001 N003 2
R3 N002 N003 10
R4 N002 0 5
R5 N003 0 4

.ac dec 10 10 10k
.end