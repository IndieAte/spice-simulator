* Basic Test Circuit

V1 N001 0 5
R1 N001 N002 100k
R2 N002 0 300k
R3 N001 N003 1k
Q1 N003 N002 N004 PNP
R4 N004 0 2k

.ac dec 20 10 10k
.end
