* Basic Test Circuit

V1 N001 0 AC(1 0)
V2 N002 N001 3
D1 N002 N003 diode
R1 N003 0 5k

.ac dec 5 1 20
.model diode D (Is=1n)
.end