* Basic Test Circuit

V1 N001 N002 AC(2 0)
R1 N001 0 100
R2 N002 0 200

.ac dec 20 10 1k
.end