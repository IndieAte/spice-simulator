* Test Circuit

V1 N001 0 1
V2 N04 2
R1 N001 N002 0 1
R2 N003 2
MOSFET N002 N004 N003

.ac dec 5 1 20
.end