* Test Circuit

V1 N001 0 2
V2 N004 0 3
R1 N001 N002 10
M1 N002 N004 0 NMOS

.ac dec 5 1 20
.end